module RF(
    input         clk, 
    input         rst,
    input         RFWr,                // 写信号
    input  [4:0]  A1, A2, A3, reg_sel, // 读寄存器号
    input  [31:0] WD,                  // 写寄存器值
    output [31:0] RD1, RD2, reg_data   // 读寄存器值
);

    reg [31:0] rf[31:0];
    integer i;

    always @(posedge clk, posedge rst)
        if (rst) begin    //  reset
            for (i=1; i<32; i=i+1) rf[i] <= 0;
        end
        else if (RFWr && A3 != 0) begin
            rf[A3] <= WD;
            // $display("r[00-07]=0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X", rf[0], rf[1], rf[2], rf[3], rf[4], rf[5], rf[6], rf[7]);
            // $display("r[08-15]=0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X", rf[8], rf[9], rf[10], rf[11], rf[12], rf[13], rf[14], rf[15]);
            // $display("r[16-23]=0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X", rf[16], rf[17], rf[18], rf[19], rf[20], rf[21], rf[22], rf[23]);
            // $display("r[24-31]=0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X, 0x%8X", rf[24], rf[25], rf[26], rf[27], rf[28], rf[29], rf[30], rf[31]);
            $display("r[%2d] = 0x%8X,", A3, WD); // 仿真时调试用，显示寄存器修改情况
        end
    

    assign RD1 = (A1 != 0) ? rf[A1] : 0;
    assign RD2 = (A2 != 0) ? rf[A2] : 0;
    assign reg_data = (reg_sel != 0) ? rf[reg_sel] : 0; // 下板 debug 用
endmodule 
